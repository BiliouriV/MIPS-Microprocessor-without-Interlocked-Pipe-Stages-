library verilog;
use verilog.vl_types.all;
entity control_bypass_ex is
    port(
        bypassA         : out    vl_logic_vector(1 downto 0);
        bypassB         : out    vl_logic_vector(1 downto 0);
        idex_rs         : in     vl_logic_vector(4 downto 0);
        idex_rt         : in     vl_logic_vector(4 downto 0);
        exmem_rd        : in     vl_logic_vector(4 downto 0);
        memwb_rd        : in     vl_logic_vector(4 downto 0);
        exmem_regwrite  : in     vl_logic;
        memwb_regwrite  : in     vl_logic
    );
end control_bypass_ex;
